module main #()();

  
endmodule
