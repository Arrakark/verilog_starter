`timescale 10ns/100ps
module main_tb;



endmodule
